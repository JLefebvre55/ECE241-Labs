module hex_decoder(c, display);
    input [3:0] c;
    output [6:0] display;
    // 3j0 2h1 1g2 0f3
    assign display[0] = ~(
        (~c[3] & ~c[2] & ~c[1] & ~c[0]) | //0
        // (~c[3] & ~c[2] & ~c[1] &  c[0]) | //1
        (~c[3] & ~c[2] &  c[1] & ~c[0]) | //2
        (~c[3] & ~c[2] &  c[1] &  c[0]) | //3
        // (~c[3] &  c[2] & ~c[1] & ~c[0]) | //4
        (~c[3] &  c[2] & ~c[1] &  c[0]) | //5
        (~c[3] &  c[2] &  c[1] & ~c[0]) | //6
        (~c[3] &  c[2] &  c[1] &  c[0]) | //7
        ( c[3] & ~c[2] & ~c[1] & ~c[0]) | //8
        ( c[3] & ~c[2] & ~c[1] &  c[0]) | //9
        ( c[3] & ~c[2] &  c[1] & ~c[0]) | //A
        // ( c[3] & ~c[2] &  c[1] &  c[0]) | //B
        ( c[3] &  c[2] & ~c[1] & ~c[0]) | //C
        // ( c[3] &  c[2] & ~c[1] &  c[0]) | //D
        ( c[3] &  c[2] &  c[1] & ~c[0]) | //E
        ( c[3] &  c[2] &  c[1] &  c[0])   //F
    );
    assign display[1] = ~(
        (~c[3] & ~c[2] & ~c[1] & ~c[0]) | //0
        (~c[3] & ~c[2] & ~c[1] &  c[0]) | //1
        (~c[3] & ~c[2] &  c[1] & ~c[0]) | //2
        (~c[3] & ~c[2] &  c[1] &  c[0]) | //3
        (~c[3] &  c[2] & ~c[1] & ~c[0]) | //4
        // (~c[3] &  c[2] & ~c[1] &  c[0]) | //5
        // (~c[3] &  c[2] &  c[1] & ~c[0]) | //6
        (~c[3] &  c[2] &  c[1] &  c[0]) | //7
        ( c[3] & ~c[2] & ~c[1] & ~c[0]) | //8
        ( c[3] & ~c[2] & ~c[1] &  c[0]) | //9
        ( c[3] & ~c[2] &  c[1] & ~c[0]) | //A
        // ( c[3] & ~c[2] &  c[1] &  c[0]) | //B
        // ( c[3] &  c[2] & ~c[1] & ~c[0]) | //C
        ( c[3] &  c[2] & ~c[1] &  c[0])   //D
        // ( c[3] &  c[2] &  c[1] & ~c[0]) | //E
        // ( c[3] &  c[2] &  c[1] &  c[0])   //F
    );
    assign display[2] = ~(
        (~c[3] & ~c[2] & ~c[1] & ~c[0]) | //0
        (~c[3] & ~c[2] & ~c[1] &  c[0]) | //1
        // (~c[3] & ~c[2] &  c[1] & ~c[0]) | //2
        (~c[3] & ~c[2] &  c[1] &  c[0]) | //3
        (~c[3] &  c[2] & ~c[1] & ~c[0]) | //4
        (~c[3] &  c[2] & ~c[1] &  c[0]) | //5
        (~c[3] &  c[2] &  c[1] & ~c[0]) | //6
        (~c[3] &  c[2] &  c[1] &  c[0]) | //7
        ( c[3] & ~c[2] & ~c[1] & ~c[0]) | //8
        ( c[3] & ~c[2] & ~c[1] &  c[0]) | //9
        ( c[3] & ~c[2] &  c[1] & ~c[0]) | //A
        ( c[3] & ~c[2] &  c[1] &  c[0]) | //B
        // ( c[3] &  c[2] & ~c[1] & ~c[0]) | //C
        ( c[3] &  c[2] & ~c[1] &  c[0])   //D
        // ( c[3] &  c[2] &  c[1] & ~c[0]) | //E
        // ( c[3] &  c[2] &  c[1] &  c[0])   //F
    );
    assign display[3] = ~(
        (~c[3] & ~c[2] & ~c[1] & ~c[0]) | //0
        // (~c[3] & ~c[2] & ~c[1] &  c[0]) | //1
        (~c[3] & ~c[2] &  c[1] & ~c[0]) | //2
        (~c[3] & ~c[2] &  c[1] &  c[0]) | //3
        // (~c[3] &  c[2] & ~c[1] & ~c[0]) | //4
        (~c[3] &  c[2] & ~c[1] &  c[0]) | //5
        (~c[3] &  c[2] &  c[1] & ~c[0]) | //6
        // (~c[3] &  c[2] &  c[1] &  c[0]) | //7
        ( c[3] & ~c[2] & ~c[1] & ~c[0]) | //8
        ( c[3] & ~c[2] & ~c[1] &  c[0]) | //9
        // ( c[3] & ~c[2] &  c[1] & ~c[0]) | //A
        ( c[3] & ~c[2] &  c[1] &  c[0]) | //B
        ( c[3] &  c[2] & ~c[1] & ~c[0]) | //C
        ( c[3] &  c[2] & ~c[1] &  c[0]) | //D
        ( c[3] &  c[2] &  c[1] & ~c[0])   //E
        // ( c[3] &  c[2] &  c[1] &  c[0])   //F
    );
    assign display[4] = ~(
        (~c[3] & ~c[2] & ~c[1] & ~c[0]) | //0
        // (~c[3] & ~c[2] & ~c[1] &  c[0]) | //1
        (~c[3] & ~c[2] &  c[1] & ~c[0]) | //2
        // (~c[3] & ~c[2] &  c[1] &  c[0]) | //3
        // (~c[3] &  c[2] & ~c[1] & ~c[0]) | //4
        // (~c[3] &  c[2] & ~c[1] &  c[0]) | //5
        (~c[3] &  c[2] &  c[1] & ~c[0]) | //6
        // (~c[3] &  c[2] &  c[1] &  c[0]) | //7
        ( c[3] & ~c[2] & ~c[1] & ~c[0]) | //8
        // ( c[3] & ~c[2] & ~c[1] &  c[0]) | //9
        ( c[3] & ~c[2] &  c[1] & ~c[0]) | //A
        ( c[3] & ~c[2] &  c[1] &  c[0]) | //B
        ( c[3] &  c[2] & ~c[1] & ~c[0]) | //C
        ( c[3] &  c[2] & ~c[1] &  c[0]) | //D
        ( c[3] &  c[2] &  c[1] & ~c[0]) | //E
        ( c[3] &  c[2] &  c[1] &  c[0])   //F
    );
    assign display[5] = ~(
        (~c[3] & ~c[2] & ~c[1] & ~c[0]) | //0
        // (~c[3] & ~c[2] & ~c[1] &  c[0]) | //1
        // (~c[3] & ~c[2] &  c[1] & ~c[0]) | //2
        // (~c[3] & ~c[2] &  c[1] &  c[0]) | //3
        (~c[3] &  c[2] & ~c[1] & ~c[0]) | //4
        (~c[3] &  c[2] & ~c[1] &  c[0]) | //5
        (~c[3] &  c[2] &  c[1] & ~c[0]) | //6
        // (~c[3] &  c[2] &  c[1] &  c[0]) | //7
        ( c[3] & ~c[2] & ~c[1] & ~c[0]) | //8
        ( c[3] & ~c[2] & ~c[1] &  c[0]) | //9
        ( c[3] & ~c[2] &  c[1] & ~c[0]) | //A
        ( c[3] & ~c[2] &  c[1] &  c[0]) | //B
        ( c[3] &  c[2] & ~c[1] & ~c[0]) | //C
        // ( c[3] &  c[2] & ~c[1] &  c[0]) | //D
        ( c[3] &  c[2] &  c[1] & ~c[0]) | //E
        ( c[3] &  c[2] &  c[1] &  c[0])   //F
    );
    assign display[6] = ~(
        // (~c[3] & ~c[2] & ~c[1] & ~c[0]) | //0
        // (~c[3] & ~c[2] & ~c[1] &  c[0]) | //1
        (~c[3] & ~c[2] &  c[1] & ~c[0]) | //2
        (~c[3] & ~c[2] &  c[1] &  c[0]) | //3
        (~c[3] &  c[2] & ~c[1] & ~c[0]) | //4
        (~c[3] &  c[2] & ~c[1] &  c[0]) | //5
        (~c[3] &  c[2] &  c[1] & ~c[0]) | //6
        // (~c[3] &  c[2] &  c[1] &  c[0]) | //7
        ( c[3] & ~c[2] & ~c[1] & ~c[0]) | //8
        ( c[3] & ~c[2] & ~c[1] &  c[0]) | //9
        ( c[3] & ~c[2] &  c[1] & ~c[0]) | //A
        ( c[3] & ~c[2] &  c[1] &  c[0]) | //B
        // ( c[3] &  c[2] & ~c[1] & ~c[0]) | //C
        ( c[3] &  c[2] & ~c[1] &  c[0]) | //D
        ( c[3] &  c[2] &  c[1] & ~c[0]) | //E
        ( c[3] &  c[2] &  c[1] &  c[0])   //F
    );
    
endmodule